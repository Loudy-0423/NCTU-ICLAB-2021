//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//      (C) Copyright NCTU OASIS Lab      
//            All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   2021 ICLAB fall Course Online Test
//   Author    : Echin-Wang    (echinwang861025@gmail.com)
//               ShaoWen-Cheng (shaowen0213@gmail.com)
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`ifdef RTL
	`timescale 1ns/10ps
	`include "GF.v"
	`define CYCLE_TIME 10.0
`endif
`ifdef GATE
	`timescale 1ns/10ps
	`include "GF_SYN.v"
	`define CYCLE_TIME 10.0
`endif

module PATTERN(
   clk,
   rst_n,
   in_valid,
   in_x,
   in_y,
   out_valid,
   out_x,
   out_y,
   out_area
     
);

output reg clk,rst_n,in_valid;
output reg [9:0] in_x,in_y;
input out_valid;
input [24:0] out_area;
input [9:0] out_x,out_y;

//================================================================
// wires & registers
//================================================================

reg [9:0] golden_x,golden_y;
reg [20:0] golden_area;
reg [2:0] golden_cycle;


//================================================================
// parameters & integer
//================================================================

integer total_cycles;
integer patcount;
integer cycles;
integer a, b, c, i, k, input_file,output_file;
integer gap;

parameter PATNUM=2000;
//================================================================
// clock
//================================================================
always	#(`CYCLE_TIME/2.0) clk = ~clk;
initial	clk = 0;
//================================================================
// initial
//================================================================
initial begin
	rst_n    = 1'b1;
	in_valid = 1'b0;
	in_x     =  'dx;
	in_y     =  'dx;
	
	force clk = 0;
	total_cycles = 0;
	reset_task;
	input_file=$fopen("../00_TESTBED/in_2000.txt","r");
  	output_file=$fopen("../00_TESTBED/out_2000.txt","r");
    @(negedge clk);
	
	for (patcount=0;patcount<PATNUM;patcount=patcount+1) begin
		input_data;
		wait_out_valid;
		check_ans;
		$display("\033[0;36mPASS PATTERN NO.%4d,\033[m \033[1;32m Cycles: %3d\033[m", patcount ,cycles);
	end
	#(1000);
	YOU_PASS_task;
	$finish;
end

task reset_task ; begin
	#(10); rst_n = 0;

	#(10);
	if((out_x !== 0) || (out_y !== 0) || (out_valid !== 0) ) begin
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                                        FAIL!                                                               ");
		$display ("                                                  Output signal should be 0 after initial RESET at %8t                                      ",$time);
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                        MMMMMMWKdc:::::::cclxOkl:::::::::::cokxl:;,,;:lxOxol:::::::::::cc:::::::::::co0WMMWKxl::::cokXWMMMMM                ");
		$display ("                        MMMMMM0,  ..........    ...........     ......      ...........  ............ ,0WO:.  .....  .oKMMMM                ");
		$display ("                        MMMMMMO. ,OXXK000KK0o.  cKXK000000k,  ;x0KKKK0x;   .oXXK000000x..o00KXXXK000c .xx. .lO0OkO0x;. ;KMMM                ");
		$display ("                        MMMMMMk. ;KMO;...;kWWd. oWWd'......  ;KMKc''cOXO;  .xMNo'......  ...,kWNd'... ,d;  ckx;..'xWNc .dWMM                ");
		$display ("                        MMMMMMk. ;KM0:,,,cOWNl  oWWx;,,,,,.  'kWNkoc::;'.  .xMNd,,,,,'.     .dWNc .,co0Xl.      .;OWK: .dWMM                ");
		$display ("                        MMMMMMk. ;KMNKKNWWKx;.  lWWX000000l.  .:dk0XNNKd'  .xMWX00000O:  .. .dWNc '0MMMMNOo:.  ;kNKd' .lXMMM                ");
		$display ("                        MMMMMMk. ;KMO,.c0WXo.   lWWd......   'cc. ..,dNMk. .xMXl......   .. .dWNc '0MMMMMMMO' 'ONk' .;kNMMMM                ");
		$display ("                        MMMMMMk. ;KMk.  'kWWO,  oWWd'....... lNWOc'';xNWx. .xMXl.......     .dWNc '0MMMMMMMO. .ox:  ;KMMMMMM                ");
		$display ("                        MMMMMMO. ,0Nd.   .oKXO,.cXNK0000000c  ;x0XKKKKOl.  .oXXK000000O;    .oXK: ,0MMMMMMMO. ,OXl  ;XMMMMMM                ");
		$display ("                        MMMMMM0,  ...  ',  .... ............    ......      ...........  ..  .... :XMMMMMMMK,  ...  lNMMMMMM                ");
		$display ("                        MMMMMMWKoc:::cdXXkl:::::::::::::::::lxxo:;,,;:cdkxlc:::::::::::coO0dc:::cxXMMMMMMMMWKoc:::cxXMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWMMMMMMMWWWWWMMMMMMMMMMMMWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0xdxOKKKKXXNNNNNWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNxcccclllllooooooddxkOO0XWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXOolccccccccc::;,',;:::::cxXWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKkdlc::ccc:cc:::;;;;::;,;:,,cxKWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0xddl::ccccccc::::::::::;;::'',lONMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKdodolcclllollc::::::::::::c:'.',ckNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNx;coololc:;:::::::::::::;,,;,..',;ckNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXd;:c:::;;,'.';lodoolcccc:,,,''',,;;cOWMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0c,,,,,,:looddxkO00Oxdlcc:;;;;;;;;;;;l0WMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXx:''',;:coddxOO00KKK0Okdolc:::::::::::;cxXWMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMWO:'..';clooododxOO000K00Okxdoccc::::c:;;;;;lkXWMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMWO,.....;lolllc::ldkOOOOOOkkxdolc::;;::;;;;;;::lxKNMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMW0:....':lllc;'.,coxOOOOOkkxdoolc:;;;;,,;;;;:::::lxKWMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMWXxl;;;::;;,,,;coxkO0OOOkxdoolc::;;;,,,;;:::::::::lOXWMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWNXKOoc::cloxkOOOOOOkxdollc:;;;,,,,;;:::::::::::cdKWMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0doodxkkkOOOkkxxdolc:;;;;;,,;;;:::::::::;,,;:l0WMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKkxxxkkkkkxxxddolc::;;;;;;;;:::ccc:::::;,,,,,,l0WMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKkkkkkkkkkxxddoolc::::;:::ccccccccccc:;,,,,,',;lKWMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNKOkkkkkkOOkkxddoollcccllllooooollcc:;,',,,,,',;:xNMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKOkkkkkOO0OOkxxdddooodddxddddoollc;;,,,,,,'',;::l0WMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKOOkkkkOO00OOkkxxxxxxkkkxxddoolcc:;;;;;,''',;;::;oKWMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKOOkkkkOOOOOOOkkkkkkkkxxddooollccc::;;;,..,;;:::;;dNMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNKOOOOOOOOOOOOOOOkkkkxxddddoooooolc::;;,''',;::;;,';kWMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMN0kkOOOOOkkOOOOOOkkkkkkxxxxdxxxddlc:;;,,'',;;;;;,'..:0MMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMN0kkkkkkOOOOOkkkkkkkkkOkkkkkxkxxoc:;;;,,',,;;;;,''..'dNMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMN0kkxxxxkOOOOkOOOOOkkkkkkkkkkxxoc::;;,,,,,;;;;,,'''',oXMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0xxdddxkkkkkkOOOkkkkkkkkkkkxdoc:;;;;,,,,;;;;,,''',,,lKMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKxoooodxkkkkkkkkxxxxxxxkxxxdoc::;;;,,,,;;;;,,,,',,,,:0MMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKdoooooddxkkxxxxdxxdddxxdoolc:;;;;,,,,,;;;;,,,,,,,,,lKMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKdodddddddxxxxxxxddddddoolc:::;;;;,,,,;;;;;,,,,,,,,;dNMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0ooddxxxdddddddxxxxxddoolc::::;;;,,'',,;;;,,,,,,''';OWMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0dddxxxxxdooooooddddddollc:::;;;,'.'',,,,,'',,,,,,;dXMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0ddxxkkkxoc:cllooooooodolcc:::;,'...'''''''',,,;,:xNMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0ddxxkkkdc;'':ccllllclodolcc::;;,.....''''',,,,,:kNMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWNKOkddxxkkxo:,''',;clllllodolccc:;;,.....''''','',cOWMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMWWNXKOkxolllodxxxkdc;,'''',:llllloddolcc:;;,.....'''''',:xXWMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMWX0Okxdocc::cldxxxxxoc,'',;:clloooodddolc::;;,......''.';dKWMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMW0oll:cloddxOK0xxdddoc:;;cloooooddddddollc:;;;,.......':xKWMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMWKxxxod0XNWMMNOdddooc:;:coodddxxxxxxddolc:;,,,'....';lOXWMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMWMMWMMMMWNXOddddoc:;:loxxxxxxxxxxdddolc:;,,,...;oOXWMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMWWWNXKOkxdoodddoooccoxkOOkkkkxxdlloolcc:,,,;:oOXWMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMWXkxkxdolclloddddx0XXXXNNNNNNXXXK0kdoolc:;,,lONWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMNd;:oooooodxxxxxOXWMMMMMMMMMMMMMMMMXkolc:,,lKWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMWOoooddddxxxxkOKWMMMMMMMMMMMMMMMMMMNkolc:;:OWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMWKxodddodddkKNMMMMMMMMMMMMMMMMMMMMXkolc:;:OWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMWXOkkxdxk0NWMMMMMMMMMMMMMMMMMMMMMKdolc:;:kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWWMMMMMMMMMMMMMMMMMMMMMMMW0dol:;,:OWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNOdolc;,oXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKkddoc::kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKxdddoc:l0MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXdoddocclxNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");
		$display ("                        MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXoccll:oKNWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM                ");

		#(100);
	    $finish ;
	end
	
	#(10); rst_n = 1 ;
	#(3.0); release clk;
end endtask

task input_data ; 
	begin
		gap = $urandom_range(1,5);
		repeat(gap)@(negedge clk);
		in_valid = 'b1;
		for(i=0;i<6;i=i+1)begin
			a = $fscanf(input_file,"%d %d",in_x,in_y);
			@(negedge clk);
		end
		in_valid     = 'b0;
		in_x         = 'bx;
		in_y         = 'bx;
	end 
endtask

task wait_out_valid ; 
begin
	cycles = 0;
	while(out_valid === 0)begin
		cycles = cycles + 1;
		if(cycles == 10000) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                                                                                            ");
			$display ("                                                     The execution latency are over 10000 cycles                                              ");
			$display ("                                                                                                                                            ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end
	@(negedge clk);
	end
	total_cycles = total_cycles + cycles;
end 
endtask

task check_ans ; 
begin
	golden_cycle = 1;
	b = $fscanf(output_file,"%d",golden_area);
	if(out_valid === 1 && out_area !== golden_area) begin
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                        FAIL!                                                               ");
			$display ("                                                                   Pattern NO.%03d                                                     ", patcount);
			$display ("                                                       Your output -> area: %d                               ", out_area);
			$display ("                                                     Golden output -> area: %d                                ", golden_area);
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXX0kolccldkKXX0xolccldOKXXXXXXXXXXXXXXXXKkollokOdllldO0xolccldO0kolllloxkdlllooolllllllldOXXXXXXXX0xollodOKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXOc'.';;;,..,l:..';;;,..;xKXXXXXXXXXXXXXKo..,'... .;.....';;;,.....',;,....';;. .,;;;;;;'.,kXXXXXOc'.,;;,'.;xKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXx'.:O0kxx0Ko. .cOKkxk00o..oKXXXXXXXXXXXXKc :XO'   oNd. :OKOxx00d. :0XWNo. :XWWd.:XXkdddd:..xXXXXO;.;kOolk0o..xXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXX0; cN0;   'lo' lN0;...,OWd..xXXXXXXXXXXXXKc :XKl,';kWd.:XXc....xNk.:0NNN0;.kNNWd.:NKc,,,'. ,OXXXXk' .,. .oXO'.oXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXk'.xWx. .oxkk:.xWx..o, oWO..dXXXXXXXXXXXXKc :XNOxxkKWd.oWO..l: :NK;:0NKkKkdKOOWd.:NNOxxxd, :0XXXXKkl;. ;O0o'.:0XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXX0; cXK:..'lKWd.lNK:...,OWd..xXXXXXXXXXXXXKc :X0'  .dWx.:XXl...'xNk.:0N0ckNW0cxWd.:NO'      ,OXXXXXXXd..ok, 'dKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXx'.:k0kxk0Kk; .cO0Oxk00l..lKXXXXXXXXXXXXKc ;XO'   oNd. ;kKOxk00d. :0XO':XNo.oNd.:XXkddddl..oXXXXXXXd..dx' cKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXOc...,;,,...;;..',;,'..;xKXXXXXXXXXXXXXKo..,'... .,. ....,;,'.....',' .',. .,. .,;;;;;;'..xXXXXXXXk'.''..oKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXX0xoccclox0XXOxlcccldOKXXXXXXXXXXXXXXXXKxlllokOdllldO0xocccldk0xlllllllllllllllllllllllokKXXXXXXXKkolllxKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKK0000000000000KKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKK00OkxdoolllllccccccccccllllodxkO0KXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK0kdolc:cloddxkO0KXXXXXXXXXXXXXK0Okdolcclox0KXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKkolcloxO00KNWWMMMMMMMMMMMMMMMMMMMMMMMMWNX0Odc:cd0XXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKxlclx0NWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXOdlclkKXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKOl:o0WMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWNOoclkKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKx:cONMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNOc:d0XXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0o:oKWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKo;l0XXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0o;xNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXo;o0XXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKx:oXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNd;dKXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKXKKKKKKKKKKKKKKKKKKKKKKKKKKKXKKKKKKKKKKKKKKKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXk:lKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM0::kXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXX0kdolllllllllllllllllllllllllllllllllllllllllllllllloox0XXXXXXXXXXXXXXXXXXXXXXXXXXXXOc;kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNd;dKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXKOdccdkO000000000000000000000000000000000000000000000O00d:o0XXXXXXXXXXXXXXXXXXXXXXXXXXXk:cKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM0clKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXX0o:cd0NWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMMMXl;xKXXXXXXXXXXXXXXXXXXXXXXXXXKd;dNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXo:OXXXXXXXXXXXXX");
			$display ("XXXXXXXXXKd;,codddddddddddddddddddddddddddddddddddddddddddddolxXMMMNd,lKXXXXXXXXXXXXXXXXXXXXXXXXXOc:0MMMMMMMMMMMMMWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNx:xXXXXXXXXXXXXX");
			$display ("XXXXXXXXXKdckKKKKKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKKKKKOl',kWMMM0:c0XXXXXXXXXXXXXXXXXXXXXXXXXk;cKWMMMMMMMMWXXNNNNNOxKWMMMMMWWWNXXK000OkONMMMMMMMMMMMMMMMMMMMMMMWx:dKXXXXXXXXXXXX");
			$display ("XXXXXXXXXKdc0MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXd;,,lXMMMXo:xXXXXXXXXXXXXXXXXXXXXXXXXXx;,ldxkOOO000xcdKNWMWO:;ldddxdooooooollllc:dXMMMMMMMMMMMMMMMMMMMMMWx:xXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXxckWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXd:oOoc0MMMWO:l0XXXXXXXXXXXXXXXXXXXXXXXXk;,oxoloollc;;l0WMMMMWO:':dkO000KXXNNNWWNXd:kWMMMMMMMMMMMMMMMMMMMMXo:kXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXkcdNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKo:kNWOcxWMMMNo:xXXXXXXXXXXXXXXXXXXXXXXXX0l;xOldXWWN0clKMMMMMMMWx:xX0KWMMMMMMMMMMWXd:kWMMMMMMMMMMMMMMMMMMMWk:lKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXX0c;odddddddddddddddxkkkkkkkkOOO0000000KKKKK00kc:kWMMXocKMMMWk;oKXXXXXXXXXXXXXXXXXXXXXXXXx:o0O0NWWXd:kWMMMMMMMM0c:kKNWMMMMMMMMWNOlcxNMMMMMMMMMMMMMMMMMMMMKl;xXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXKx;,okOOOOOkkkkxxxxxxkxxxxxxxxddoollllooooollc,cKMMMWk:dNMMWO:l0XXXXXXXXXXXXXXXXXXXXXXXXO:,cllooolokXWMMMMMMMMWOc:okOKXXK0OxdollxKNMMMMMMMMMMMMMMMMMMMMNd;o0XXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXX0l;xNMMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWWWWWWWWWXocOWMMM0:lXMMMNo:xXXXXXXXXXXXXXXXXXXXXXXXX0o,ckOOO0XNMMMMMMMMMMMMWXOxoooooolloxOKNWMMMMMMMMMMMMMMMMMMMMMXd:o0XXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXk:cKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWOcoNMMMNoc0MMMWOcoKXXXXXXXXXXXXXXXXXXXXXXXX0lcOWMMMMMMMMMMWWWWWMMMMMMWWNNNNNWWMMMMMMMMMMMMMMMMMMMMMMMMWXo;l0XXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXKo;kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMKccKMMMWOcdNMMMXo:kXXXXXXXXXXXXXXXXXXXXXXXXXOcc0WMMMWK0OOkkxxxxkkOXWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0l:d0XXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXx;oNMMMMMMMMWWWWWWWWWMMMMMMMMMMMMMMMMMWMMMMNx:xNMMMNdcOWMMWx;oKXXXXXXXXXXXXXXXXXXXXXXXXKx:oXWWXd;,''',,,,'''';lx0NMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXkccxKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXX0l:OWMMMMMW0ooooooooddxddxkkkkkkkOKX0xxKMMMMKccKMMMWO:dNMMWO::OXXXXXXXXXXXXXXXXXXXXXXXXXKx:lkxlldxdxkO00Okxdoolc:oOXWMMMMMMMMMMMMMMMMMMMMMMMMW0l:oOXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXx:oNMMMMMNd;o0K0000OOOkkxkkkkkkkk0k;.;0MMMMNx:xNMMM0c:0MMMXo:kXXXXXXXXXXXXXXXXXXXXXXXXXXKx;'':0WMMWKkddddx0NWWN0o:l0NMMMMMMMMMMMMMMMMMMMMMW0ocoOKXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXX0l:0WMMMMXo:0MMMMMMMMMMMMMMMMMMMMNd;,;xWMMMM0::0WMMNd:kWMMWk:dKXXXXXXXXXXXXXXXXXXXXXXXXXXKo,.:0WMMWXOkxxxdkNMMMMN0o:dXWMMMMMMMMMMMMMMMMMN0o:lOKXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXKd;oXMMMMKclKMMMMMMMMMMMMMMMMMMMMKl:oclKMMMMXo;kWMMMKclXMMMXlcOXXXXXXXXXXXXXXXXXXXXXXXXXX0l;c:cdKWMMMMMMMMMMMMMMMWNkcl0WMMMMMMMMMMMMMWXkl;;dKXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXOccKMMMWk:xNMMMMMMMMMMMMMMMMMMMM0:c0x:kWMMMWO:oNMMMNd:kWMMWk:oKXXXXXXXXXXXXXXXXXXXXXXXXXk:cO0dccoONWMMMMMMMMMMMMMMW0l:kNMMMMMMMMWNKOdc,'.:OXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXKd:xWMMNoc0MMMMMMMMMMMMMMMMMMMMWO:dNO:dNMMMMXo:OWMMW0clXMMMKccOXXXXXXXXXXXXXXXXXXXXXXXXXx;l0XXKkocld0XWMMMMMMMMMMMMWXx:oKWMMWX0xllcldxd:';xXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXOccKWM0clXMMMMMMMMMMMMMMMMMMMMWkckWO:dNMMMMW0clXMMMNo;kWMMXl;xXXXXXXXXXXXXXXXXXXXXXXXXKo,oKXXXXK0xollodOKXNWWWWWWWWWXd;cxxdl:;;lxOKXXXOc,l0XXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXKd:dNWO;oNMMMMMMMMMMMMMMMMMMMMWxl0Nx:OWMMMMMNo:OWMMWk;oNMMWx;oKXXXXXXXXXXXXXXXXXXXXXXXKo;dKXXXXXXXXKkdlllllolloooolllc;'''.';oOKXXXXXXKd,,dKXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXO::0Nd;xWMMMMMMMMMMMMMMMMMMMMXllKKllKMMMMMMWx;oNMMMKllKMMMKl:OXXXXXXXXXXXXXXXXXXXXXXXKl:kXXXXXXXXXXXXXXK0OOkxxkkxxkkkkxl,':kKXXXXXXXXKd,';dKXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXX0l;kXo:OMMMMMMMMMMMMMMMMMMMMM0cdNk:xWMMMMMMMXlcKMMMWx:xNMMWx:dKXXXXXXXXXXXXXXXXXXXXXX0c:kXXXXXXXXXXXXXXXXXXXXXXXXXXXXKkc,,l0XXXXXXXXXKo;:;;xXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXk:okclKMMMMMMMMMMMMMMMMMMMMWxcONxcOMMMMMMMMWkcxWMMMXlc0MMM0ccOXXXXXXXXXXXXXXXXXXXXXXO:cOXXXXXXXXXXXXXXXXXXXXXXXXXXXOo:cdl;dKXXXXXXXXO:ckx:ckXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXKo::;dNMMMMMMMMMMMMMMMMMMMMNocKXl:OMMMMMMMMMXllKMMMWx;xWMMNo;dKXXXXXXXXXXXXXXXXXXXXXO:l0XXXXXXXXXXXXXXXXXXXXXXXXKOdccxKX0l:xKXXXXXXKx;oKKx;cOXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXk:':OWMMMMMMMMMMMMMMMMMMMMKcoXXc:0MMMMMMMMMWk:xNMMWO:oNMMWx;oKXXXXXXXXXXXXXXXXXXXXXO:l0XXXXXXXXXXXXXXXXXXXXXXX0d:cxKXXXXk::kXXXXXXKo;xXX0c,dKXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXX0l'cKMMMMMMMMMMMMMMMMMMMMMO;oX0:oNMMMMMMMMMM0clXMMMXoc0WMMKcc0XXXXXXXXXXXXXXXXXXXXXO:cOXXXXXXXXXXXXXXXXXXXXK0dccx0XXXXXXKd;oKXXXXXOc:OXXXx;cOXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKo,oNMMMMMMMMMMMMMMMMMMMMWx;dKd:OWMMMMMMMMMMNdc0MMMWOcdNMWKlcOXXXXXXXXXXXXXXXXXXXXX0l:kXXXXXXXXXXXXXXXXXXXOo:cx0XXXXXXXXX0l:xXXXXXk;l0XXXKo:xXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKl;xWMMMMMMMMMMMMMMMMMMMMNo;kKlcKMMMMMMMMMMMM0coKWMMXo:OXklcxKXXXXXXXXXXXXXXXXXXXXXKo;dKXXXXXXXXXXXXXXXKOoclx0XXXXXXXXXXXXk:cOXXXKo,l0XXXXk:lKXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKo;kWMMMMMMMMMMMMMMMMMMMMNoc0O:lOKKKKKKKKKKKKOl,;ldxxl,:ccd0XXXXXXXXXXXXXXXXXXXXXXXKo,oKXXXXXXXXXXXXXKkl:cx0XXXXXXXXXXXXXX0l;dKXX0c;xKXXXX0l:kXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXX0lc0MMMMMMMMMMMMMMMMMMMMMKloKd,',;;;,;;;;;;;;,,'''''',;lx0XXXXXXXXXXXXXXXXXXXXXXXXXXd;l0XXXXXXXXXXX0xlclkKXXXXXXXXXXXXXXXXKd,c0XKd:o0XXXXXKo;dKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXk:lXMMMMMMMMMMMMMMMMMMMMWOcx0c,lxxxxxxxxxxxxxxxxxxxxxkOKKXXKKKK000OO00KKXXXXXXXXXXXXk;c0XXXXXXXXKOoccdOKXXXXXXXXXXXXXXXXXXXOc:OXOccOXXXXXXKo,oKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXKd:xWMMMMMMMMMMMMMMMMMMMMWx:dx;':cccccccccccccccloooooooooooooollc:;:ccllloxO0KXXXXXXOc:OXXXXXX0xlcok0XXXXXXXXXXXXXXXXXXXXXXKd:xOc;dKXXXXXXKd;oKXXXXXXXXXXXXXXXXXX");
			$display ("XKKKKKKKKKKKKKKKKKOc;d00KKKXXXXXXXXXXKKKKKK0o,;:;;;;;;;;;;;;;;;;cdk0KKKXKKKKKXXXXXK0lcOXK0Okdl:ckXXXXXXKo;oKXX0koccdOKXXXXXXXXXXXXXXXXXXXXXXXXXx:lo;cOXXXXKXXKd;cOXKKKKKKKKKKKKKKKXX");
			$display ("dooolllllooooooolc;;coddddxxxkkkkkxxxxxxxxxxkxlo0KXXXKXKKKKKKKKXNKdxXWMMMMMMMMMMMMMNocKMMMWWWKc,cooddddoc,;lol:,,:loddddddddddddddddddddddddddoc,,,,:odoolllll:,;clllllllllcccccccco");
			$display ("KKKKKKKKKKKKKKK0o;cONWWWMWWWWWWWMWWWWWWWWWWWMXooXMMMMMMMMMMMMMMMMNkccxOO0000000000Okc;oddddddo::lxkOOOOOOkkOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOkxdodkOOOOOOOOOOOOOOkkxxolc:,'',,;;:;;");
			$display ("MMMMMMMMMMMMMMNx:l0NNNWWWWNNNNXKKKKKKKKKKKKKK0l:lddxxxxxxxxxxxxxxxdl:codxkkkkkkkkkkkxxxxxxxxkOKXWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWMMMMWNNXKOOkxdddooodddxxxkO0KXXNx:");
			$display ("MMMMMMMMMMMMMW0ocoxxdddxxxddddoollooddoooooddxxxxxxkOOOOOOOkkkkkOO0KXNWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWNXK0kxddddooloodxxxxkO0XNWWWMMMMMMMMMWk:");
			$display ("MMMMMMMMMMMMMMWNNNNNXXXXXXNNNNNNNNWWWWWWWWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWNXK0OkkxdoooooooodxkOO0XNWWMMMMMMMMMMMMMMMMMMMMMWk:");
			$display ("MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWX0dc,'',;lxO0XNWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWk:");
			@(negedge clk);
			$finish;
	end
    while(out_valid === 1) begin
		
		c = $fscanf(output_file,"%d %d",golden_x,golden_y);
		if(	(out_x !== golden_x) || (out_y !== golden_y)) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                        FAIL!                                                               ");
			$display ("                                                                   Pattern NO.%03d                                                     ", patcount);
			$display ("                                                       Your output -> out_x: %d,  out_y: %d                                ", out_x, out_y);
			$display ("                                                     Golden output -> out_x: %d,  out_y: %d                                ", golden_x, golden_y);
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXX0kolccldkKXX0xolccldOKXXXXXXXXXXXXXXXXKkollokOdllldO0xolccldO0kolllloxkdlllooolllllllldOXXXXXXXX0xollodOKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXOc'.';;;,..,l:..';;;,..;xKXXXXXXXXXXXXXKo..,'... .;.....';;;,.....',;,....';;. .,;;;;;;'.,kXXXXXOc'.,;;,'.;xKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXx'.:O0kxx0Ko. .cOKkxk00o..oKXXXXXXXXXXXXKc :XO'   oNd. :OKOxx00d. :0XWNo. :XWWd.:XXkdddd:..xXXXXO;.;kOolk0o..xXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXX0; cN0;   'lo' lN0;...,OWd..xXXXXXXXXXXXXKc :XKl,';kWd.:XXc....xNk.:0NNN0;.kNNWd.:NKc,,,'. ,OXXXXk' .,. .oXO'.oXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXk'.xWx. .oxkk:.xWx..o, oWO..dXXXXXXXXXXXXKc :XNOxxkKWd.oWO..l: :NK;:0NKkKkdKOOWd.:NNOxxxd, :0XXXXKkl;. ;O0o'.:0XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXX0; cXK:..'lKWd.lNK:...,OWd..xXXXXXXXXXXXXKc :X0'  .dWx.:XXl...'xNk.:0N0ckNW0cxWd.:NO'      ,OXXXXXXXd..ok, 'dKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXx'.:k0kxk0Kk; .cO0Oxk00l..lKXXXXXXXXXXXXKc ;XO'   oNd. ;kKOxk00d. :0XO':XNo.oNd.:XXkddddl..oXXXXXXXd..dx' cKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXOc...,;,,...;;..',;,'..;xKXXXXXXXXXXXXXKo..,'... .,. ....,;,'.....',' .',. .,. .,;;;;;;'..xXXXXXXXk'.''..oKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXX0xoccclox0XXOxlcccldOKXXXXXXXXXXXXXXXXKxlllokOdllldO0xocccldk0xlllllllllllllllllllllllokKXXXXXXXKkolllxKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKK0000000000000KKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKK00OkxdoolllllccccccccccllllodxkO0KXXXXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK0kdolc:cloddxkO0KXXXXXXXXXXXXXK0Okdolcclox0KXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKkolcloxO00KNWWMMMMMMMMMMMMMMMMMMMMMMMMWNX0Odc:cd0XXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKxlclx0NWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXOdlclkKXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKOl:o0WMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWNOoclkKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKx:cONMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNOc:d0XXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0o:oKWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKo;l0XXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX0o;xNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXo;o0XXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKx:oXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNd;dKXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKXKKKKKKKKKKKKKKKKKKKKKKKKKKKXKKKKKKKKKKKKKKKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXk:lKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM0::kXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXX0kdolllllllllllllllllllllllllllllllllllllllllllllllloox0XXXXXXXXXXXXXXXXXXXXXXXXXXXXOc;kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNd;dKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXKOdccdkO000000000000000000000000000000000000000000000O00d:o0XXXXXXXXXXXXXXXXXXXXXXXXXXXk:cKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM0clKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXX0o:cd0NWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMMMXl;xKXXXXXXXXXXXXXXXXXXXXXXXXXKd;dNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXo:OXXXXXXXXXXXXX");
			$display ("XXXXXXXXXKd;,codddddddddddddddddddddddddddddddddddddddddddddolxXMMMNd,lKXXXXXXXXXXXXXXXXXXXXXXXXXOc:0MMMMMMMMMMMMMWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNx:xXXXXXXXXXXXXX");
			$display ("XXXXXXXXXKdckKKKKKKXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXKKKKKOl',kWMMM0:c0XXXXXXXXXXXXXXXXXXXXXXXXXk;cKWMMMMMMMMWXXNNNNNOxKWMMMMMWWWNXXK000OkONMMMMMMMMMMMMMMMMMMMMMMWx:dKXXXXXXXXXXXX");
			$display ("XXXXXXXXXKdc0MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXd;,,lXMMMXo:xXXXXXXXXXXXXXXXXXXXXXXXXXx;,ldxkOOO000xcdKNWMWO:;ldddxdooooooollllc:dXMMMMMMMMMMMMMMMMMMMMMWx:xXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXxckWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXd:oOoc0MMMWO:l0XXXXXXXXXXXXXXXXXXXXXXXXk;,oxoloollc;;l0WMMMMWO:':dkO000KXXNNNWWNXd:kWMMMMMMMMMMMMMMMMMMMMXo:kXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXkcdNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKo:kNWOcxWMMMNo:xXXXXXXXXXXXXXXXXXXXXXXXX0l;xOldXWWN0clKMMMMMMMWx:xX0KWMMMMMMMMMMWXd:kWMMMMMMMMMMMMMMMMMMMWk:lKXXXXXXXXXXXXX");
			$display ("XXXXXXXXXX0c;odddddddddddddddxkkkkkkkkOOO0000000KKKKK00kc:kWMMXocKMMMWk;oKXXXXXXXXXXXXXXXXXXXXXXXXx:o0O0NWWXd:kWMMMMMMMM0c:kKNWMMMMMMMMWNOlcxNMMMMMMMMMMMMMMMMMMMMKl;xXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXKx;,okOOOOOkkkkxxxxxxkxxxxxxxxddoollllooooollc,cKMMMWk:dNMMWO:l0XXXXXXXXXXXXXXXXXXXXXXXXO:,cllooolokXWMMMMMMMMWOc:okOKXXK0OxdollxKNMMMMMMMMMMMMMMMMMMMMNd;o0XXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXX0l;xNMMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWWWWWWWWWXocOWMMM0:lXMMMNo:xXXXXXXXXXXXXXXXXXXXXXXXX0o,ckOOO0XNMMMMMMMMMMMMWXOxoooooolloxOKNWMMMMMMMMMMMMMMMMMMMMMXd:o0XXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXk:cKMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWOcoNMMMNoc0MMMWOcoKXXXXXXXXXXXXXXXXXXXXXXXX0lcOWMMMMMMMMMMWWWWWMMMMMMWWNNNNNWWMMMMMMMMMMMMMMMMMMMMMMMMWXo;l0XXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXKo;kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMKccKMMMWOcdNMMMXo:kXXXXXXXXXXXXXXXXXXXXXXXXXOcc0WMMMWK0OOkkxxxxkkOXWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0l:d0XXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXx;oNMMMMMMMMWWWWWWWWWMMMMMMMMMMMMMMMMMWMMMMNx:xNMMMNdcOWMMWx;oKXXXXXXXXXXXXXXXXXXXXXXXXKx:oXWWXd;,''',,,,'''';lx0NMMMMMMMMMMMMMMMMMMMMMMMMMMMMWXkccxKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXX0l:OWMMMMMW0ooooooooddxddxkkkkkkkOKX0xxKMMMMKccKMMMWO:dNMMWO::OXXXXXXXXXXXXXXXXXXXXXXXXXKx:lkxlldxdxkO00Okxdoolc:oOXWMMMMMMMMMMMMMMMMMMMMMMMMW0l:oOXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXx:oNMMMMMNd;o0K0000OOOkkxkkkkkkkk0k;.;0MMMMNx:xNMMM0c:0MMMXo:kXXXXXXXXXXXXXXXXXXXXXXXXXXKx;'':0WMMWKkddddx0NWWN0o:l0NMMMMMMMMMMMMMMMMMMMMMW0ocoOKXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXX0l:0WMMMMXo:0MMMMMMMMMMMMMMMMMMMMNd;,;xWMMMM0::0WMMNd:kWMMWk:dKXXXXXXXXXXXXXXXXXXXXXXXXXXKo,.:0WMMWXOkxxxdkNMMMMN0o:dXWMMMMMMMMMMMMMMMMMN0o:lOKXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXKd;oXMMMMKclKMMMMMMMMMMMMMMMMMMMMKl:oclKMMMMXo;kWMMMKclXMMMXlcOXXXXXXXXXXXXXXXXXXXXXXXXXX0l;c:cdKWMMMMMMMMMMMMMMMWNkcl0WMMMMMMMMMMMMMWXkl;;dKXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXOccKMMMWk:xNMMMMMMMMMMMMMMMMMMMM0:c0x:kWMMMWO:oNMMMNd:kWMMWk:oKXXXXXXXXXXXXXXXXXXXXXXXXXk:cO0dccoONWMMMMMMMMMMMMMMW0l:kNMMMMMMMMWNKOdc,'.:OXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXKd:xWMMNoc0MMMMMMMMMMMMMMMMMMMMWO:dNO:dNMMMMXo:OWMMW0clXMMMKccOXXXXXXXXXXXXXXXXXXXXXXXXXx;l0XXKkocld0XWMMMMMMMMMMMMWXx:oKWMMWX0xllcldxd:';xXXXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXOccKWM0clXMMMMMMMMMMMMMMMMMMMMWkckWO:dNMMMMW0clXMMMNo;kWMMXl;xXXXXXXXXXXXXXXXXXXXXXXXXKo,oKXXXXK0xollodOKXNWWWWWWWWWXd;cxxdl:;;lxOKXXXOc,l0XXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXKd:dNWO;oNMMMMMMMMMMMMMMMMMMMMWxl0Nx:OWMMMMMNo:OWMMWk;oNMMWx;oKXXXXXXXXXXXXXXXXXXXXXXXKo;dKXXXXXXXXKkdlllllolloooolllc;'''.';oOKXXXXXXKd,,dKXXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXO::0Nd;xWMMMMMMMMMMMMMMMMMMMMXllKKllKMMMMMMWx;oNMMMKllKMMMKl:OXXXXXXXXXXXXXXXXXXXXXXXKl:kXXXXXXXXXXXXXXK0OOkxxkkxxkkkkxl,':kKXXXXXXXXKd,';dKXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXX0l;kXo:OMMMMMMMMMMMMMMMMMMMMM0cdNk:xWMMMMMMMXlcKMMMWx:xNMMWx:dKXXXXXXXXXXXXXXXXXXXXXX0c:kXXXXXXXXXXXXXXXXXXXXXXXXXXXXKkc,,l0XXXXXXXXXKo;:;;xXXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXk:okclKMMMMMMMMMMMMMMMMMMMMWxcONxcOMMMMMMMMWkcxWMMMXlc0MMM0ccOXXXXXXXXXXXXXXXXXXXXXXO:cOXXXXXXXXXXXXXXXXXXXXXXXXXXXOo:cdl;dKXXXXXXXXO:ckx:ckXXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXKo::;dNMMMMMMMMMMMMMMMMMMMMNocKXl:OMMMMMMMMMXllKMMMWx;xWMMNo;dKXXXXXXXXXXXXXXXXXXXXXO:l0XXXXXXXXXXXXXXXXXXXXXXXXKOdccxKX0l:xKXXXXXXKx;oKKx;cOXXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXk:':OWMMMMMMMMMMMMMMMMMMMMKcoXXc:0MMMMMMMMMWk:xNMMWO:oNMMWx;oKXXXXXXXXXXXXXXXXXXXXXO:l0XXXXXXXXXXXXXXXXXXXXXXX0d:cxKXXXXk::kXXXXXXKo;xXX0c,dKXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXX0l'cKMMMMMMMMMMMMMMMMMMMMMO;oX0:oNMMMMMMMMMM0clXMMMXoc0WMMKcc0XXXXXXXXXXXXXXXXXXXXXO:cOXXXXXXXXXXXXXXXXXXXXK0dccx0XXXXXXKd;oKXXXXXOc:OXXXx;cOXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKo,oNMMMMMMMMMMMMMMMMMMMMWx;dKd:OWMMMMMMMMMMNdc0MMMWOcdNMWKlcOXXXXXXXXXXXXXXXXXXXXX0l:kXXXXXXXXXXXXXXXXXXXOo:cx0XXXXXXXXX0l:xXXXXXk;l0XXXKo:xXXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKl;xWMMMMMMMMMMMMMMMMMMMMNo;kKlcKMMMMMMMMMMMM0coKWMMXo:OXklcxKXXXXXXXXXXXXXXXXXXXXXKo;dKXXXXXXXXXXXXXXXKOoclx0XXXXXXXXXXXXk:cOXXXKo,l0XXXXk:lKXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXKo;kWMMMMMMMMMMMMMMMMMMMMNoc0O:lOKKKKKKKKKKKKOl,;ldxxl,:ccd0XXXXXXXXXXXXXXXXXXXXXXXKo,oKXXXXXXXXXXXXXKkl:cx0XXXXXXXXXXXXXX0l;dKXX0c;xKXXXX0l:kXXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXX0lc0MMMMMMMMMMMMMMMMMMMMMKloKd,',;;;,;;;;;;;;,,'''''',;lx0XXXXXXXXXXXXXXXXXXXXXXXXXXd;l0XXXXXXXXXXX0xlclkKXXXXXXXXXXXXXXXXKd,c0XKd:o0XXXXXKo;dKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXXk:lXMMMMMMMMMMMMMMMMMMMMWOcx0c,lxxxxxxxxxxxxxxxxxxxxxkOKKXXKKKK000OO00KKXXXXXXXXXXXXk;c0XXXXXXXXKOoccdOKXXXXXXXXXXXXXXXXXXXOc:OXOccOXXXXXXKo,oKXXXXXXXXXXXXXXXXXX");
			$display ("XXXXXXXXXXXXXXXXXXKd:xWMMMMMMMMMMMMMMMMMMMMWx:dx;':cccccccccccccccloooooooooooooollc:;:ccllloxO0KXXXXXXOc:OXXXXXX0xlcok0XXXXXXXXXXXXXXXXXXXXXXKd:xOc;dKXXXXXXKd;oKXXXXXXXXXXXXXXXXXX");
			$display ("XKKKKKKKKKKKKKKKKKOc;d00KKKXXXXXXXXXXKKKKKK0o,;:;;;;;;;;;;;;;;;;cdk0KKKXKKKKKXXXXXK0lcOXK0Okdl:ckXXXXXXKo;oKXX0koccdOKXXXXXXXXXXXXXXXXXXXXXXXXXx:lo;cOXXXXKXXKd;cOXKKKKKKKKKKKKKKKXX");
			$display ("dooolllllooooooolc;;coddddxxxkkkkkxxxxxxxxxxkxlo0KXXXKXKKKKKKKKXNKdxXWMMMMMMMMMMMMMNocKMMMWWWKc,cooddddoc,;lol:,,:loddddddddddddddddddddddddddoc,,,,:odoolllll:,;clllllllllcccccccco");
			$display ("KKKKKKKKKKKKKKK0o;cONWWWMWWWWWWWMWWWWWWWWWWWMXooXMMMMMMMMMMMMMMMMNkccxOO0000000000Okc;oddddddo::lxkOOOOOOkkOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOkxdodkOOOOOOOOOOOOOOkkxxolc:,'',,;;:;;");
			$display ("MMMMMMMMMMMMMMNx:l0NNNWWWWNNNNXKKKKKKKKKKKKKK0l:lddxxxxxxxxxxxxxxxdl:codxkkkkkkkkkkkxxxxxxxxkOKXWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWMMMMWNNXKOOkxdddooodddxxxkO0KXXNx:");
			$display ("MMMMMMMMMMMMMW0ocoxxdddxxxddddoollooddoooooddxxxxxxkOOOOOOOkkkkkOO0KXNWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWWNXK0kxddddooloodxxxxkO0XNWWWMMMMMMMMMWk:");
			$display ("MMMMMMMMMMMMMMWNNNNNXXXXXXNNNNNNNNWWWWWWWWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWNXK0OkkxdoooooooodxkOO0XNWWMMMMMMMMMMMMMMMMMMMMMWk:");
			$display ("MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWX0dc,'',;lxO0XNWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWk:");
			@(negedge clk);
			$finish;
		end
		
		@(negedge clk);
		golden_cycle=golden_cycle+1;
    end
	if(golden_cycle !== 6+1) begin
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                                        FAIL!                                                               ");
		$display ("                                                                   Pattern NO.%03d                                                     ", patcount);
		$display ("	                                                         Output cycle should be 6 cycle                                              ");
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		@(negedge clk);
		$finish;
	end
end 
endtask

task YOU_PASS_task;
	begin
	$display ("WWWWWWWWWWWWWWWWWWWMMWWWWWWWWWWWWWWWWWWWWWWMMMWWWWMMMMMMMMWWWWWWWWWWNNNNNNXXXXXXKK0KNMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMWWWWN");
	$display ("WWWWWWWWWWWWWWWWWWWWWWWWWWWWWNNNNXXXXKKKK0000OOkkkkxxxddddooollllcc:::;;;,,,,'''''.;OWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMWWWWWWWWWWWWWWWWMMWMMWWWMWWWWN");
	$display ("WWWWWWWWWWWWWWWNkooolllccc:::;;;,,,,'''............................................'kWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMWWWWWWWWWN");
	$display ("WWWWWWWWWWWWWWWKc...................................................'''',,,,;;,.....xWMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWN");
	$display ("WWWWWMMWWWMMWWMXc............''',,,;;::::ccclllooodddxxxxkkkOOO000KKKXXXNNNNNNKc....dWMMWWWWWWWWWWWWWWWMMWMWWWWWWWWWWWWWWWMMWWWWWWWWWWWWMMWWWWWWWWWWWW");
	$display ("WWWWWWMWWMMMWMMNl....:kO000KKKXXXNNNNWWWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNl....oNMWWWWWWWWWWWWWWWWMWWWWWWWWWWWWWWWWWWWMMMMMWWWWWWWWMWWWWWWWWWWWWN");
	$display ("WWWWWWWMMMMWWMMNo....oNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNo....oNMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMWWMWWWWWWWWWWWWWWWWWWWWN");
	$display ("WWWWWWWWWWMWWMMNd....lNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWd....lXWWMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWMMWWWWx....cXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWx....cXWWWMMMWWMMWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMWWWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWk'...cXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWk'...:0XXXXXXNNWWWWMMWWWWWWWWWWWWWWWWWWWWWWWMMWWWWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWMWMMWk'...:KMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWk'....;c:::::ccclodxOKNWWWWWWWWWWWWWWWWWWWWMMWWWMMWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWMMWMWO,...;KMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMO,....:llooollllc::;;::ldkKNWWWWWWWWWWWWWWWMWWWWWWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWMMWWW0,...,0MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM0,....,:;;;;;:lloooooolc;;:cdONWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWMMWWW0;...,OMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMK;...'dK00Oxdlc:;;cloooooolc;;:o0NWWWWWWWWWWWWWWWWWWWWWWMWWWWWWWWWWWWWW");
	$display ("WWWWWWWWMMWWWWWMK:...'kMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMK:...'kWMMMMMMWXOdc;;:loooooolc;;cxKWWWWWWWWWWWWWWWWWWWWWWWMWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMXc....kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXc....xWMMMMMMMMMMWKxl;;coooooool:;;o0NWWWWWWWWWWWWWWWWWWWMMMWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMXc....xWMMMWNNNNWWMMMMMMMMMWNNWMMMMMMMMMWNNNWMMMMMMMMWNNNNWMMMMXl....dWMMMMMMMMMMMMMWKd:;:loooooooc;;lONWMWWMWWMMWWWWWWWMWWWWWWWWWWWWN");
	$display ("WWWWWWWWWWWWWWWMNl....dWMKl,,,,;;;cxXMMMMKo;,,;xNMMMMXxc;;;;;ckNMMNOl;;;;;:ldXMNo....dWMMMMMMMMMMMMMMMWXkc,:loooooool;;l0NWMMWWMWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMNo....oNMx.,xkddxxc.:KMMXc.:kx,.dWMMX:.cxxxkx;.cXNo.;xkxxkc,.;0No....oNMMMMMMMMMMMMMMMMMMNkc,:looooollc;,l0WWWWWWWWWWWWWWWWWWWWWWMWWWW");
	$display ("WWWWWWWWWWWWWWWMNd....lNMx.:NO,.:0N:.xMNo.:KXXO'.kWMk.,KXo,:ol..OK,.kNx;;ooc'.dNd....lNMMMMMMMMMMMMMMMMMMMMNx:,cool;'..',';dXWWWWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWx....lXMx.:NKdoxKk''OWk.,0K:oXk.,0WO..:xOkkx:..OK; ,dkOkxl;..dNx....;OXWMMMMMMMMMMMMMMMMMMMWKo,;l:..   ..'':kNWWMMWWMWWWMMWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWk'...cXMx.:N0l::;,:OW0,.kN0xkXNd.:Ko.'l;..:0Nc.ox..c:..,kNWd.:Xk'...'llcokKWMMMMMMMMMMMMMMMMMNk;,;..   ...',,lKWWWWWWWWWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMWk'...:KMx.:Kx.'dOKWMX:.oKd''',kKc.lx''k0xox0k,.k0;.o0kdd00x:.oNO'...'cc..:ood0NMMMMMMMMMMMMMMMW0c''.. .;:..;:,:OWWWMWWWMWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMWO,...;KMO,.,'.oWMMMMK:.',.;kx,.,'.lXOc,;:::;,:OWWKl,,:::;,';xNMO,....lxd:co;.'cxKWMMMMMMMMMMMMMWXl''..    .'cl;,xNWWMMWMWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMW0,...;0MWXOOOKWMMMMMMX0OO0NMMX0OO0NMMWX0kkkOXWMMMMWX0kkkOKXNMMM0,...'d00kdodc,:l:l0WMMMMMMMMMMMMMXl',,.. ..,lol:,dXMWMMWWWWWWWWWWWWWW");
	$display ("WWWWWWWMMWWWWWMMW0;...,OMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMK;...'o000000kocl;.,o0WMMMMMMMMMMMMXl,:c:;;:loooo:,oXMMMWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWMMWWWWWWK:...'kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMK:....;llx00000OOo;cc;oXMMMMMMMMMMMMXc,coooooooooo:,oNWWMWWWWMWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWKc....kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXc....;oc;colcok0Ool:..cOWMMMMMMMMMMMK:,loooooooooo:,dNWWWWWWWWWWWWWWW");
	$display ("WWWWWWWMMWWWWWWWWXc....xWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXc....;oo;.'cc;:oookx:;;;xNMMMMMMMMMMWO;,loooooooooo:,dNWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWXl....dWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNl....dNWXKkdo;.'c::dxo:..oNMMMMMMMMMMWx,:ooooooooool;;OWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWNo....oNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNo....oNMMMMMWXOxo:';k0d,''oNMMMMMMMMMMXl'cooooooooooolOWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWNd....lNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWd....lNMMMMMMMMMWKxlccolc;,dNMMMMMMMMMM0:,loooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWWx....lXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWx....cXMMMMMMMMMMMMWKxlclxl;kWMMMMMMMMMWx,:oooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWMWx'...cXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWx....:XMMMMMMMMMMMMMMMN0dc:':0MMMMMMMMMMXl'cooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWMWk'...:KMMMMMMMMMMMMMMMMMMMMW0xx0NMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMk'...:KMMMMMMMMMMMMMMMMMWXx;'dWMMMMMMMMMMO,;ooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWMWO,...;KMMMMMMMMMMMMMMMMMMMXo,;;,oXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMO,...;0MMMMMMMMMMMMMMMMMMMMN0KWMMMMMMMMMMNl'coooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWW0,...,0MMMMMMMMMMMMMMMMMMXl':oo:,dNMMMMMMMMMMMMMMMMMMMMMMMMMMMM0,...,0MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWO,';;;;;;;:oKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWMMMMWW0;...,OMMMMMMMMMMMMMMMMMNo':oooo;;OWMMMMMMMMMMMMMMMMMMMMMMMMMMM0;...,OMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNl.,::::::cdKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWMMWMK:...'kMMMMMMMMMMMMMMMMWk,;oooool;lXMMMMMMMMMMMMMMMMMMMMMMMMMMMK:...'kWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMO,;looollldKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWMWMXc....xWMMMMMMMMMMMMMMM0;'looooooc;xWMMMMMMMMMMMMMMMMMMMWWWWWWW0:....xWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMXc.,;,,,,,cOWWWWWWWWMMWWWN");
	$display ("WWWWWWWWWWWWWWWMWWXc....xWMMMMMMMWWWWWWWXl':oooooooo;;xOOOkkkxxxdddooolllcccc:::;,.....dNWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMWx',lllllldKWWWWWWWWMMWWWN");
	$display ("WWWMMWWWWWWWWWWMWWNl....;odooolllccc:::;,.'looooooool'.......................    ......,ccclllooooddxxkO0KXNWWMMMMMMMMMMMMMMMK:':ccc::l0WMWWWWWWWWWWWN");
	$display ("WWWWMMWWWWWWWWWMMMNo.................... .;oooooooooo:. ..................... .;::cccccccccccccc::::;;;;;::cllodkOKNWMMMMMMMMWd.',;,,;:OWMWWWWWWWWWWWN");
	$display ("WWWWWMMWWWWWWWWMMMWd...............'''''..cooooooooool'.:ddddxxxkkOOOO000KKKd.'looooooooooooooooooooooooooollc::;;:clodk0XWMMM0;;loooodKWWWWWWWWWWWWWW");
	$display ("WWWWWMMWWWWWWWWWWWWKxxxkkkkOOOO0000KKXX0:.cooooooooooo:,dNMMMMMMMMMMMMMMMMMMNx:,;cloooooooooooooooooooooooooooooooolc:;;;:cok0Kl.,;,,,:OWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWMMWWWWWWMWWMMMWWWWWWWWWWWWWWWWXc.coooooooooool,;0MMMMMMMMMMMMMMMMMMMMNOl:,,:looooooooooooooooooooooooooooooooooolc:;;:,..;:cco0WWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWMWWWMMMMWWMMWWWWWWWWWWWWWWWWWNd':oooooooooooo:'dWMMMMMMMMMMMMMMMMMMMMMMN0xl:;;cloooooooooooooooooooooooooooooooooooolc;,,,,;l0WWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWMMWWMMWWWWWWWWWWWWWWWWWWWWWWWW0:,loooooooooool,:KMMMMMMMMMMMMMMMMMMMMMMMMMWXOdc;;clooooooooooooooooooooooooooooooooooooool:;c0WWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWMMWWMWWWWWWWWWWWWWWWWWWWWWWWWWNO:;looooooooooo:,xWMMMMMMMMMMMMMMMMMMMMMMMMMMMMWKxc;;cooooooooooooooooooooooooooooooooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWMMMWWWWWWWWWMWWWWWWWWWWWWWWWWWWWKo;;coooooooool,lXMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMN0d:;:loooooooooooooooooooooooooooooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWN0dc;;cloooooo;;OMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMNkc;;looooooooooooooooooooooooooooooooooxKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMWN0xl:;:loooc,oNMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMW0l;;coooooooooooooooooooooooooooooooodKWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMWWWWMMWWMMWWWWKkdkO00OkONWWWMMMMMMMMMMMMMMMMMMWWWWMMMMMMMMMMMMWKxxO0000000000000000000000000000000KNWWWWWWWWWWWWWW");
	$display ("WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMMMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWWWWWW");
	$display ("\033[1;36m----------------------------------*****************************************************----------------------------------------------\033[m");
	$display ("                                           \033[1;35m       Congratulations! \033[m               						            ");
	$display ("                                           \033[1;35mYou have passed all patterns! \033[m         						            ");
	$display ("                                           \033[0;38mYour execution cycles = %5d cycles \033[m  						            ", total_cycles);
	$display ("                                           \033[0;38mYour clock period  = %.1f ns \033[m       					                ", `CYCLE_TIME);
	$display ("                                           \033[0;38mYour total latency = %.1f ns \033[m        						            ", total_cycles*`CYCLE_TIME);
	$display ("\033[1;36m----------------------------------*****************************************************----------------------------------------------\033[m");
	
	$finish;

	end
endtask

endmodule