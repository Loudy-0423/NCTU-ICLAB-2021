
`ifdef RTL
	`timescale 1ns/10ps
	`include "MAZE.v"
    `define CYCLE_TIME 10.0
`endif
`ifdef GATE
	`timescale 1ns/10ps
	`include "MAZE_SYN.v"
    `define CYCLE_TIME 10.0
`endif

module PATTERN(
    // Output signals
	clk,
    rst_n,
	in_valid,
	in,
    // Input signals
    out_valid,
    out
);

output reg clk, rst_n, in_valid, in;
input out_valid;
input [1:0] out;

//================================================================
// wires & registers
//================================================================
reg [8:0] loc;
reg golden[288:0];

//================================================================
// parameters & integer
//================================================================

integer total_cycles;
integer patcount;
integer cycles;
integer a, b, i, k, input_file,output_file;
integer gap;

parameter PATNUM=300;//104;

//================================================================
// clock
//================================================================
always	#(`CYCLE_TIME/2.0) clk = ~clk;
initial	clk = 0;
//================================================================
// initial
//================================================================

initial begin
	rst_n    = 1'b1;
	in_valid = 1'b0;
	in     =  'dx;
	
	force clk = 0;
	total_cycles = 0;
	loc = 0;
	reset_task;
	
	
	input_file=$fopen("../00_TESTBED/input.txt","r");
  	output_file=$fopen("../00_TESTBED/input.txt","r");
    @(negedge clk);

	for (patcount=0;patcount<PATNUM;patcount=patcount+1) begin
		input_data;
		wait_out_valid;
		check_ans;
		$display("\033[0;34mPASS PATTERN NO.%4d \033[m \033[0;32m \033[m", patcount);
	end
	#(100000);//1000
	YOU_PASS_task;
	$finish;
end

task reset_task ; begin
	#(10); rst_n = 0;

	#(10);
	if((out_valid !== 0) || (out !== 0)) begin
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                                        SPEC 3 IS FAIL!                                                     ");
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		
		#(100);
	    $finish ;
	end
	
	#(10); rst_n = 1 ;
	#(3.0); release clk;
end endtask



task input_data ; 
	begin
		gap = $urandom_range(1,5);
		repeat(gap)@(negedge clk);
		in_valid = 'b1;
		for(i=0;i<289;i=i+1)begin
			/* if(out !== 0) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 4 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				repeat(2)@(negedge clk);
				$finish;
			end */
			if(out_valid === 1) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 5 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				repeat(2)@(negedge clk);
				$finish;
			end
			a = $fscanf(input_file,"%d",in);
			b = $fscanf(output_file,"%d",golden[i]);
			@(negedge clk);
		end
			
		//@(negedge clk);
		in_valid = 'b0;
		in = 'bx;
	end 
endtask





task wait_out_valid ; 
begin
	cycles = 0;
	while(out_valid === 0)begin
		cycles = cycles + 1;
		if(out !== 0) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 4 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end
		if(cycles == 3000) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 6 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end
	@(negedge clk);
	end
	//total_cycles = total_cycles + cycles;
end 
endtask



task check_ans ; 
begin
	//cycles = 0;
    while(out_valid === 1) begin
		cycles = cycles + 1;
		if(out === 0) begin
			if(golden[loc+1] === 0 || (loc+1)%17 === 0) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 7 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				@(negedge clk);
				$finish;
			end
			else begin
				loc = loc+1;
			end
		end
		else if(out === 1) begin
			if(golden[loc+17] === 0 || loc > 271) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 7 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				@(negedge clk);
				$finish;
			end
			else begin
				loc = loc+17;
			end
		end
		else if(out === 2) begin
			if(golden[loc-1] === 0 || loc%17 === 0) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 7 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				@(negedge clk);
				$finish;
			end
			else begin
				loc = loc-1;
			end
		end
		else if(out === 3) begin
			if(golden[loc-17] === 0 || loc < 17) begin
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				$display ("                                                                   SPEC 7 IS FAIL!                                                          ");
				$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
				@(negedge clk);
				$finish;
			end
			else begin
				loc = loc-17;
			end
		end
		
		if(/* total_cycles +  */cycles == 3000) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 6 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end

	@(negedge clk);
    end
	if(out_valid === 0) begin
		cycles = cycles + 1;
		if(out !== 0) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 4 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end
		if(loc !== 288) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 7 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			@(negedge clk);
			$finish;
		end
		if(/* total_cycles +  */cycles == 3000) begin
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                                   SPEC 6 IS FAIL!                                                          ");
			$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2)@(negedge clk);
			$finish;
		end
	end
	//total_cycles = total_cycles + cycles;
	loc = 0;
end 
endtask






task YOU_PASS_task;
	begin
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$display ("                                                  Congratulations!                						            ");
	$display ("                                           You have passed all patterns!          						            ");
	$display ("----------------------------------------------------------------------------------------------------------------------");
	$finish;

	end
endtask


endmodule